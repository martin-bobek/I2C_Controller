library ieee;
use ieee.std_logic_1164.all;

entity application is
  port (
    clk     : in std_logic;
    buttons : in std_logic_vector(1 downto 0)
  );
end;

architecture rtl of application is
begin

end;